BZh91AY&SY9To= j_�Py��g�����P��@��5=ORmI��OҞ(H4 4j 9�14L�2da0M4����sbh0�2d��`�i���!����a2dɑ��4�# C ��M Гʟ�4�OP�@��oI/đԋr�P�D
�?l
D�I $_�D�Z�NX5b���4�ܫ�f(�{L7��ߥ8E���g�=]wu��.qqi[��7�̙#�
#Z�ޕ��E���Z�w�;�6l9����RH�!1,{���$��0w��Q2L�d��rcT"Wd@v�ek*VB�.-�vT��b�LzA4�w:��h��ޙ5�����8���=�C���B_-5�@p�A��Z*{	v$Ҁ^�@Z�$�L�R��m�p�8z)J��Z��r��
�������X�Kf�bW��X�@k�BÏ��E��:lY�f�nb��[�ym}��@uJ���E����f���D��g�����.#�37�Gh�#\����$���J��o}�*�E������%�8��e�G��M��ć�M�"RC�y��D{=7аoG �x�3�t&e�1ί>q+*�M���ކ�B�K�eH�f����y~n�P��l0*pA�R0;v�Pw�����%�b��b>:��!��2Y�i��<VK�!�aS��)���Ha\I�8��"��Y���0�����i.X��0�!��@vD$U	IL���%%D��+)�ô�l�;F�(�S��=Wr�s.-�O� �X���:�7G��t�BB;0,kD�������o�MC]P�*fړ� ��cű[wd���/�ڰ.!2��Jp�WAyn�ׁ��Vn8�{
Ij�`~2��|Y/�w9 ����h�������I��J�L�6�������.���e�j�\Y���.�p� r��z